/home/andrey/Anna/Programming/fpga/core/pipistrello/minsoc1/minsoc/prj/../rtl/verilog/adv_debug_sys/Hardware/altera_virtual_jtag/rtl/vhdl//altera_virtual_jtag.vhd
